module our;
   initial begin $display("My first ever design."); $finish; end
endmodule
